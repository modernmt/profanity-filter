horornas	1.0
kukarnas	1.0
djävelns	1.0
fittornas	1.0
jävlarnas	1.0
kukens	1.0
snorrarna	1.0
ludrets	1.0
bögens	1.0
kukar	0.97529536
jävelns	0.9705882
horans	0.969697
kuk	0.92904806
negerns	0.9285714
kuken	0.9251935
fittorna	0.9142857
knullas	0.9113924
fitta	0.9022789
kukarna	0.8965517
jävlarna	0.89649224
jäveln	0.89558685
röv	0.88606155
fittans	0.875
fittan	0.872093
neger	0.86733
jävel	0.866652
hora	0.8658408
röven	0.86032563
knulla	0.85483587
horan	0.8479685
negern	0.84659094
horor	0.8453441
hororna	0.8358209
djäveln	0.8181818
knullande	0.8130081
djävel	0.7883212
ludret	0.7619048
muttor	0.75
jävla	0.72856236
jävlar	0.72448766
luder	0.7094017
fnask	0.68
åt helvete	0.67248416
rövar	0.65229887
blatte	0.6511628
djävla	0.6371308
mutta	0.63225806
ludren	0.6
fnasket	0.5959596
blatten	0.57894737
fnasken	0.5625
negrernas	0.5555556
bögen	0.5450237
knullandes	0.5
muttorna	0.5
muttan	0.46
balle	0.40458015
bögarna	0.4
fnaskets	0.4
bögar	0.3814774
djävlarna	0.32520324
svartskalle	0.31034482
djävlar	0.29386893
snorren	0.2857143
bög	0.24637681
blattarna	0.23529412
svartskallarna	0.23076923
ballen	0.2173913
negrer	0.19911504
rövarna	0.19565217
svartskallen	0.18181819
tattare	0.1764706
bögarnas	0.1764706
tattaren	0.16666667
ballarna	0.1594203
snorre	0.15517241
negrerna	0.14634146
snorrar	0.14285715
svartskallar	0.13636364
ballar	0.12548262
blattar	0.05
muttans	0.0
djävlarnas	0.0
tattarnas	0.0
svartskallarnas	0.0
ballarnas	0.0
ludrens	0.0
snorrarnas	0.0
tattarens	0.0
muttornas	0.0
blattarnas	0.0
snorrens	0.0
ballens	0.0
rövarnas	0.0
rövens	0.0
fnaskens	0.0
tattarna	0.0
svartskallens	0.0
blattens	0.0
